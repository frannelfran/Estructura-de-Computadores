module alu(output wire [3:0] R, output wire zero, c_out, sign, input wire [3:0] A, B, input wire c_in,
          input wire [1:0] ALUOP, input wire l);

endmodule