/* 
  3.1. Implementar un “Full-Adder” de la manera más simple posible (operador concatenación ‘{…}’), con el
  prototipo
*/

module fa(output wire c_out, sum, input wire a, b, c_in);







endmodule